module Sqrt_Finer_Lookup(
    input wire [31:0] sqrt_input,
    output logic [11:0] sqrt_output);

    always_comb begin
        if ((sqrt_input > 31'd1) && (sqrt_input <= 31'd4)) begin
                sqrt_output = 11'd1;
        end else if ((sqrt_input > 31'd4) && (sqrt_input <= 31'd9)) begin
                sqrt_output = 11'd2;
        end else if ((sqrt_input > 31'd9) && (sqrt_input <= 31'd16)) begin
                sqrt_output = 11'd3;
        end else if ((sqrt_input > 31'd16) && (sqrt_input <= 31'd25)) begin
                sqrt_output = 11'd4;
        end else if ((sqrt_input > 31'd25) && (sqrt_input <= 31'd36)) begin
                sqrt_output = 11'd5;
        end else if ((sqrt_input > 31'd36) && (sqrt_input <= 31'd49)) begin
                sqrt_output = 11'd6;
        end else if ((sqrt_input > 31'd49) && (sqrt_input <= 31'd64)) begin
                sqrt_output = 11'd7;
        end else if ((sqrt_input > 31'd64) && (sqrt_input <= 31'd81)) begin
                sqrt_output = 11'd8;
        end else if ((sqrt_input > 31'd81) && (sqrt_input <= 31'd100)) begin
                sqrt_output = 11'd9;
        end else if ((sqrt_input > 31'd100) && (sqrt_input <= 31'd121)) begin
                sqrt_output = 11'd10;
        end else if ((sqrt_input > 31'd121) && (sqrt_input <= 31'd144)) begin
                sqrt_output = 11'd11;
        end else if ((sqrt_input > 31'd144) && (sqrt_input <= 31'd169)) begin
                sqrt_output = 11'd12;
        end else if ((sqrt_input > 31'd169) && (sqrt_input <= 31'd196)) begin
                sqrt_output = 11'd13;
        end else if ((sqrt_input > 31'd196) && (sqrt_input <= 31'd225)) begin
                sqrt_output = 11'd14;
        end else if ((sqrt_input > 31'd225) && (sqrt_input <= 31'd256)) begin
                sqrt_output = 11'd15;
        end else if ((sqrt_input > 31'd256) && (sqrt_input <= 31'd289)) begin
                sqrt_output = 11'd16;
        end else if ((sqrt_input > 31'd289) && (sqrt_input <= 31'd324)) begin
                sqrt_output = 11'd17;
        end else if ((sqrt_input > 31'd324) && (sqrt_input <= 31'd361)) begin
                sqrt_output = 11'd18;
        end else if ((sqrt_input > 31'd361) && (sqrt_input <= 31'd400)) begin
                sqrt_output = 11'd19;
        end else if ((sqrt_input > 31'd400) && (sqrt_input <= 31'd441)) begin
                sqrt_output = 11'd20;
        end else if ((sqrt_input > 31'd441) && (sqrt_input <= 31'd484)) begin
                sqrt_output = 11'd21;
        end else if ((sqrt_input > 31'd484) && (sqrt_input <= 31'd529)) begin
                sqrt_output = 11'd22;
        end else if ((sqrt_input > 31'd529) && (sqrt_input <= 31'd576)) begin
                sqrt_output = 11'd23;
        end else if ((sqrt_input > 31'd576) && (sqrt_input <= 31'd625)) begin
                sqrt_output = 11'd24;
        end else if ((sqrt_input > 31'd625) && (sqrt_input <= 31'd676)) begin
                sqrt_output = 11'd25;
        end else if ((sqrt_input > 31'd676) && (sqrt_input <= 31'd729)) begin
                sqrt_output = 11'd26;
        end else if ((sqrt_input > 31'd729) && (sqrt_input <= 31'd784)) begin
                sqrt_output = 11'd27;
        end else if ((sqrt_input > 31'd784) && (sqrt_input <= 31'd841)) begin
                sqrt_output = 11'd28;
        end else if ((sqrt_input > 31'd841) && (sqrt_input <= 31'd900)) begin
                sqrt_output = 11'd29;
        end else if ((sqrt_input > 31'd900) && (sqrt_input <= 31'd961)) begin
                sqrt_output = 11'd30;
        end else if ((sqrt_input > 31'd961) && (sqrt_input <= 31'd1024)) begin
                sqrt_output = 11'd31;
        end else if ((sqrt_input > 31'd1024) && (sqrt_input <= 31'd1089)) begin
                sqrt_output = 11'd32;
        end else if ((sqrt_input > 31'd1089) && (sqrt_input <= 31'd1156)) begin
                sqrt_output = 11'd33;
        end else if ((sqrt_input > 31'd1156) && (sqrt_input <= 31'd1225)) begin
                sqrt_output = 11'd34;
        end else if ((sqrt_input > 31'd1225) && (sqrt_input <= 31'd1296)) begin
                sqrt_output = 11'd35;
        end else if ((sqrt_input > 31'd1296) && (sqrt_input <= 31'd1369)) begin
                sqrt_output = 11'd36;
        end else if ((sqrt_input > 31'd1369) && (sqrt_input <= 31'd1444)) begin
                sqrt_output = 11'd37;
        end else if ((sqrt_input > 31'd1444) && (sqrt_input <= 31'd1521)) begin
                sqrt_output = 11'd38;
        end else if ((sqrt_input > 31'd1521) && (sqrt_input <= 31'd1600)) begin
                sqrt_output = 11'd39;
        end else if ((sqrt_input > 31'd1600) && (sqrt_input <= 31'd1681)) begin
                sqrt_output = 11'd40;
        end else if ((sqrt_input > 31'd1681) && (sqrt_input <= 31'd1764)) begin
                sqrt_output = 11'd41;
        end else if ((sqrt_input > 31'd1764) && (sqrt_input <= 31'd1849)) begin
                sqrt_output = 11'd42;
        end else if ((sqrt_input > 31'd1849) && (sqrt_input <= 31'd1936)) begin
                sqrt_output = 11'd43;
        end else if ((sqrt_input > 31'd1936) && (sqrt_input <= 31'd2025)) begin
                sqrt_output = 11'd44;
        end else if ((sqrt_input > 31'd2025) && (sqrt_input <= 31'd2116)) begin
                sqrt_output = 11'd45;
        end else if ((sqrt_input > 31'd2116) && (sqrt_input <= 31'd2209)) begin
                sqrt_output = 11'd46;
        end else if ((sqrt_input > 31'd2209) && (sqrt_input <= 31'd2304)) begin
                sqrt_output = 11'd47;
        end else if ((sqrt_input > 31'd2304) && (sqrt_input <= 31'd2401)) begin
                sqrt_output = 11'd48;
        end else if ((sqrt_input > 31'd2401) && (sqrt_input <= 31'd2500)) begin
                sqrt_output = 11'd49;
        end else if ((sqrt_input > 31'd2500) && (sqrt_input <= 31'd2601)) begin
                sqrt_output = 11'd50;
        end else if ((sqrt_input > 31'd2601) && (sqrt_input <= 31'd2704)) begin
                sqrt_output = 11'd51;
        end else if ((sqrt_input > 31'd2704) && (sqrt_input <= 31'd2809)) begin
                sqrt_output = 11'd52;
        end else if ((sqrt_input > 31'd2809) && (sqrt_input <= 31'd2916)) begin
                sqrt_output = 11'd53;
        end else if ((sqrt_input > 31'd2916) && (sqrt_input <= 31'd3025)) begin
                sqrt_output = 11'd54;
        end else if ((sqrt_input > 31'd3025) && (sqrt_input <= 31'd3136)) begin
                sqrt_output = 11'd55;
        end else if ((sqrt_input > 31'd3136) && (sqrt_input <= 31'd3249)) begin
                sqrt_output = 11'd56;
        end else if ((sqrt_input > 31'd3249) && (sqrt_input <= 31'd3364)) begin
                sqrt_output = 11'd57;
        end else if ((sqrt_input > 31'd3364) && (sqrt_input <= 31'd3481)) begin
                sqrt_output = 11'd58;
        end else if ((sqrt_input > 31'd3481) && (sqrt_input <= 31'd3600)) begin
                sqrt_output = 11'd59;
        end else if ((sqrt_input > 31'd3600) && (sqrt_input <= 31'd3721)) begin
                sqrt_output = 11'd60;
        end else if ((sqrt_input > 31'd3721) && (sqrt_input <= 31'd3844)) begin
                sqrt_output = 11'd61;
        end else if ((sqrt_input > 31'd3844) && (sqrt_input <= 31'd3969)) begin
                sqrt_output = 11'd62;
        end else if ((sqrt_input > 31'd3969) && (sqrt_input <= 31'd4096)) begin
                sqrt_output = 11'd63;
        end else if ((sqrt_input > 31'd4096) && (sqrt_input <= 31'd4225)) begin
                sqrt_output = 11'd64;
        end else if ((sqrt_input > 31'd4225) && (sqrt_input <= 31'd4356)) begin
                sqrt_output = 11'd65;
        end else if ((sqrt_input > 31'd4356) && (sqrt_input <= 31'd4489)) begin
                sqrt_output = 11'd66;
        end else if ((sqrt_input > 31'd4489) && (sqrt_input <= 31'd4624)) begin
                sqrt_output = 11'd67;
        end else if ((sqrt_input > 31'd4624) && (sqrt_input <= 31'd4761)) begin
                sqrt_output = 11'd68;
        end else if ((sqrt_input > 31'd4761) && (sqrt_input <= 31'd4900)) begin
                sqrt_output = 11'd69;
        end else if ((sqrt_input > 31'd4900) && (sqrt_input <= 31'd5041)) begin
                sqrt_output = 11'd70;
        end else if ((sqrt_input > 31'd5041) && (sqrt_input <= 31'd5184)) begin
                sqrt_output = 11'd71;
        end else if ((sqrt_input > 31'd5184) && (sqrt_input <= 31'd5329)) begin
                sqrt_output = 11'd72;
        end else if ((sqrt_input > 31'd5329) && (sqrt_input <= 31'd5476)) begin
                sqrt_output = 11'd73;
        end else if ((sqrt_input > 31'd5476) && (sqrt_input <= 31'd5625)) begin
                sqrt_output = 11'd74;
        end else if ((sqrt_input > 31'd5625) && (sqrt_input <= 31'd5776)) begin
                sqrt_output = 11'd75;
        end else if ((sqrt_input > 31'd5776) && (sqrt_input <= 31'd5929)) begin
                sqrt_output = 11'd76;
        end else if ((sqrt_input > 31'd5929) && (sqrt_input <= 31'd6084)) begin
                sqrt_output = 11'd77;
        end else if ((sqrt_input > 31'd6084) && (sqrt_input <= 31'd6241)) begin
                sqrt_output = 11'd78;
        end else if ((sqrt_input > 31'd6241) && (sqrt_input <= 31'd6400)) begin
                sqrt_output = 11'd79;
        end else if ((sqrt_input > 31'd6400) && (sqrt_input <= 31'd6561)) begin
                sqrt_output = 11'd80;
        end else if ((sqrt_input > 31'd6561) && (sqrt_input <= 31'd6724)) begin
                sqrt_output = 11'd81;
        end else if ((sqrt_input > 31'd6724) && (sqrt_input <= 31'd6889)) begin
                sqrt_output = 11'd82;
        end else if ((sqrt_input > 31'd6889) && (sqrt_input <= 31'd7056)) begin
                sqrt_output = 11'd83;
        end else if ((sqrt_input > 31'd7056) && (sqrt_input <= 31'd7225)) begin
                sqrt_output = 11'd84;
        end else if ((sqrt_input > 31'd7225) && (sqrt_input <= 31'd7396)) begin
                sqrt_output = 11'd85;
        end else if ((sqrt_input > 31'd7396) && (sqrt_input <= 31'd7569)) begin
                sqrt_output = 11'd86;
        end else if ((sqrt_input > 31'd7569) && (sqrt_input <= 31'd7744)) begin
                sqrt_output = 11'd87;
        end else if ((sqrt_input > 31'd7744) && (sqrt_input <= 31'd7921)) begin
                sqrt_output = 11'd88;
        end else if ((sqrt_input > 31'd7921) && (sqrt_input <= 31'd8100)) begin
                sqrt_output = 11'd89;
        end else if ((sqrt_input > 31'd8100) && (sqrt_input <= 31'd8281)) begin
                sqrt_output = 11'd90;
        end else if ((sqrt_input > 31'd8281) && (sqrt_input <= 31'd8464)) begin
                sqrt_output = 11'd91;
        end else if ((sqrt_input > 31'd8464) && (sqrt_input <= 31'd8649)) begin
                sqrt_output = 11'd92;
        end else if ((sqrt_input > 31'd8649) && (sqrt_input <= 31'd8836)) begin
                sqrt_output = 11'd93;
        end else if ((sqrt_input > 31'd8836) && (sqrt_input <= 31'd9025)) begin
                sqrt_output = 11'd94;
        end else if ((sqrt_input > 31'd9025) && (sqrt_input <= 31'd9216)) begin
                sqrt_output = 11'd95;
        end else if ((sqrt_input > 31'd9216) && (sqrt_input <= 31'd9409)) begin
                sqrt_output = 11'd96;
        end else if ((sqrt_input > 31'd9409) && (sqrt_input <= 31'd9604)) begin
                sqrt_output = 11'd97;
        end else if ((sqrt_input > 31'd9604) && (sqrt_input <= 31'd9801)) begin
                sqrt_output = 11'd98;
        end else begin
            sqrt_output = 11'd0;
        end
    end
endmodule
