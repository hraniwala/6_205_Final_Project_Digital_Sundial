module Sqrt_Lookup(
    input wire [31:0] sqrt_input,
    output logic [31:0] sqrt_output);

    always_comb begin
        if ((sqrt_input > 32'd1000000) && (sqrt_input <= 32'd4000000)) begin
                sqrt_output = 32'd1000;
        end else if ((sqrt_input > 32'd4000000) && (sqrt_input <= 32'd9000000)) begin
                sqrt_output = 32'd2000;
        end else if ((sqrt_input > 32'd9000000) && (sqrt_input <= 32'd16000000)) begin
                sqrt_output = 32'd3000;
        end else if ((sqrt_input > 32'd16000000) && (sqrt_input <= 32'd25000000)) begin
                sqrt_output = 32'd4000;
        end else if ((sqrt_input > 32'd25000000) && (sqrt_input <= 32'd36000000)) begin
                sqrt_output = 32'd5000;
        end else if ((sqrt_input > 32'd36000000) && (sqrt_input <= 32'd49000000)) begin
                sqrt_output = 32'd6000;
        end else if ((sqrt_input > 32'd49000000) && (sqrt_input <= 32'd64000000)) begin
                sqrt_output = 32'd7000;
        end else if ((sqrt_input > 32'd64000000) && (sqrt_input <= 32'd81000000)) begin
                sqrt_output = 32'd8000;
        end else if ((sqrt_input > 32'd81000000) && (sqrt_input <= 32'd100000000)) begin
                sqrt_output = 32'd9000;
        end else if ((sqrt_input > 32'd100000000) && (sqrt_input <= 32'd121000000)) begin
                sqrt_output = 32'd10000;
        end else if ((sqrt_input > 32'd121000000) && (sqrt_input <= 32'd144000000)) begin
                sqrt_output = 32'd11000;
        end else if ((sqrt_input > 32'd144000000) && (sqrt_input <= 32'd169000000)) begin
                sqrt_output = 32'd12000;
        end else if ((sqrt_input > 32'd169000000) && (sqrt_input <= 32'd196000000)) begin
                sqrt_output = 32'd13000;
        end else if ((sqrt_input > 32'd196000000) && (sqrt_input <= 32'd225000000)) begin
                sqrt_output = 32'd14000;
        end else if ((sqrt_input > 32'd225000000) && (sqrt_input <= 32'd256000000)) begin
                sqrt_output = 32'd15000;
        end else if ((sqrt_input > 32'd256000000) && (sqrt_input <= 32'd289000000)) begin
                sqrt_output = 32'd16000;
        end else if ((sqrt_input > 32'd289000000) && (sqrt_input <= 32'd324000000)) begin
                sqrt_output = 32'd17000;
        end else if ((sqrt_input > 32'd324000000) && (sqrt_input <= 32'd361000000)) begin
                sqrt_output = 32'd18000;
        end else if ((sqrt_input > 32'd361000000) && (sqrt_input <= 32'd400000000)) begin
                sqrt_output = 32'd19000;
        end else if ((sqrt_input > 32'd400000000) && (sqrt_input <= 32'd441000000)) begin
                sqrt_output = 32'd20000;
        end else if ((sqrt_input > 32'd441000000) && (sqrt_input <= 32'd484000000)) begin
                sqrt_output = 32'd21000;
        end else if ((sqrt_input > 32'd484000000) && (sqrt_input <= 32'd529000000)) begin
                sqrt_output = 32'd22000;
        end else if ((sqrt_input > 32'd529000000) && (sqrt_input <= 32'd576000000)) begin
                sqrt_output = 32'd23000;
        end else if ((sqrt_input > 32'd576000000) && (sqrt_input <= 32'd625000000)) begin
                sqrt_output = 32'd24000;
        end else if ((sqrt_input > 32'd625000000) && (sqrt_input <= 32'd676000000)) begin
                sqrt_output = 32'd25000;
        end else if ((sqrt_input > 32'd676000000) && (sqrt_input <= 32'd729000000)) begin
                sqrt_output = 32'd26000;
        end else if ((sqrt_input > 32'd729000000) && (sqrt_input <= 32'd784000000)) begin
                sqrt_output = 32'd27000;
        end else if ((sqrt_input > 32'd784000000) && (sqrt_input <= 32'd841000000)) begin
                sqrt_output = 32'd28000;
        end else if ((sqrt_input > 32'd841000000) && (sqrt_input <= 32'd900000000)) begin
                sqrt_output = 32'd29000;
        end else if ((sqrt_input > 32'd900000000) && (sqrt_input <= 32'd961000000)) begin
                sqrt_output = 32'd30000;
        end else if ((sqrt_input > 32'd961000000) && (sqrt_input <= 32'd1024000000)) begin
                sqrt_output = 32'd31000;
        end else if ((sqrt_input > 32'd1024000000) && (sqrt_input <= 32'd1089000000)) begin
                sqrt_output = 32'd32000;
        end else if ((sqrt_input > 32'd1089000000) && (sqrt_input <= 32'd1156000000)) begin
                sqrt_output = 32'd33000;
        end else if ((sqrt_input > 32'd1156000000) && (sqrt_input <= 32'd1225000000)) begin
                sqrt_output = 32'd34000;
        end else if ((sqrt_input > 32'd1225000000) && (sqrt_input <= 32'd1296000000)) begin
                sqrt_output = 32'd35000;
        end else if ((sqrt_input > 32'd1296000000) && (sqrt_input <= 32'd1369000000)) begin
                sqrt_output = 32'd36000;
        end else if ((sqrt_input > 32'd1369000000) && (sqrt_input <= 32'd1444000000)) begin
                sqrt_output = 32'd37000;
        end else if ((sqrt_input > 32'd1444000000) && (sqrt_input <= 32'd1521000000)) begin
                sqrt_output = 32'd38000;
        end else if ((sqrt_input > 32'd1521000000) && (sqrt_input <= 32'd1600000000)) begin
                sqrt_output = 32'd39000;
        end else if ((sqrt_input > 32'd1600000000) && (sqrt_input <= 32'd1681000000)) begin
                sqrt_output = 32'd40000;
        end else if ((sqrt_input > 32'd1681000000) && (sqrt_input <= 32'd1764000000)) begin
                sqrt_output = 32'd41000;
        end else if ((sqrt_input > 32'd1764000000) && (sqrt_input <= 32'd1849000000)) begin
                sqrt_output = 32'd42000;
        end else if ((sqrt_input > 32'd1849000000) && (sqrt_input <= 32'd1936000000)) begin
                sqrt_output = 32'd43000;
        end else if ((sqrt_input > 32'd1936000000) && (sqrt_input <= 32'd2025000000)) begin
                sqrt_output = 32'd44000;
        end else if ((sqrt_input > 32'd2025000000) && (sqrt_input <= 32'd2116000000)) begin
                sqrt_output = 32'd45000;
        end else if ((sqrt_input > 32'd2116000000) && (sqrt_input <= 32'd2209000000)) begin
                sqrt_output = 32'd46000;
        end else if ((sqrt_input > 32'd2209000000) && (sqrt_input <= 32'd2304000000)) begin
                sqrt_output = 32'd47000;
        end else if ((sqrt_input > 32'd2304000000) && (sqrt_input <= 32'd2401000000)) begin
                sqrt_output = 32'd48000;
        end else if ((sqrt_input > 32'd2401000000) && (sqrt_input <= 32'd2500000000)) begin
                sqrt_output = 32'd49000;
        end else begin
            sqrt_output = 32'd0;
        end
    end
endmodule
